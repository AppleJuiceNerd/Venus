module appui

import element
