module logger

// Log severity levels
pub enum Severity as u8 {
	debug
	info
	warning
	error
	critical
}
