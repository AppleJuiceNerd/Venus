module main

import mastodon

fn main() {
	mastodon.prepare_app()
}
