module element

import src.mastodon.api
import gg
import gx
